library ieee;
use ieee.std_logic_1164.all;
--Process Al value to show on display. Display segment lights up with a 0 not 1
entity processToDisplay is

	port
	(
		al_value   : in std_logic_vector (7 downto 0);
		a0, a1 ,a2 ,a3 ,a4, a5,	a6    : out std_logic;
		b0, b1, b2, b3, b4, b5, b6    : out std_logic
		
	);

end entity;

architecture rtl of processToDisplay is

 signal rightMBs: std_logic_vector(3 downto 0);
 signal leftMBs: std_logic_vector(3 downto 0);
 
begin

	rightMBs <= al_value(3 downto 0);
	leftMBs <= al_value (7 downto 4);
	
	--for right display
	process (al_value) is
	begin
		if(rightMBs = "0000") then
			b0 <= '0';
			b1 <= '0';
			b2 <= '0';
			b3 <= '0';
			b4 <= '0';
			b5 <= '0';
			b6 <= '1';
		elsif (rightMBs = "0001") then
			b0 <= '1';
			b1 <= '0';
			b2 <= '0';
			b3 <= '1';
			b4 <= '1';
			b5 <= '1';
			b6 <= '1';
		elsif (rightMBs = "0010") then
			b0 <= '0';
			b1 <= '0';
			b2 <= '1';
			b3 <= '0';
			b4 <= '0';
			b5 <= '1';
			b6 <= '0';
		elsif (rightMBs = "0011") then
			b0 <= '0';
			b1 <= '0';
			b2 <= '0';
			b3 <= '0';
			b4 <= '1';
			b5 <= '1';
			b6 <= '0';
		elsif (rightMBs = "0100") then
			b0 <= '1';
			b1 <= '0';
			b2 <= '0';
			b3 <= '1';
			b4 <= '1';
			b5 <= '0';
			b6 <= '0';
		elsif (rightMBs = "0101") then
			b0 <= '0';
			b1 <= '1';
			b2 <= '0';
			b3 <= '0';
			b4 <= '1';
			b5 <= '0';
			b6 <= '0';
		elsif (rightMBs = "0110") then
			b0 <= '0';
			b1 <= '1';
			b2 <= '0';
			b3 <= '0';
			b4 <= '0';
			b5 <= '0';
			b6 <= '0';
		elsif (rightMBs = "0111") then
			b0 <= '0';
			b1 <= '0';
			b2 <= '0';
			b3 <= '1';
			b4 <= '1';
			b5 <= '1';
			b6 <= '1';
		elsif (rightMBs = "1000") then
			b0 <= '0';
			b1 <= '0';
			b2 <= '0';
			b3 <= '0';
			b4 <= '0';
			b5 <= '0';
			b6 <= '0';
		elsif (rightMBs = "1001") then
			b0 <= '0';
			b1 <= '0';
			b2 <= '0';
			b3 <= '1';
			b4 <= '1';
			b5 <= '0';
			b6 <= '0';
			elsif (rightMBs = "1010") then
			b0 <= '0';
			b1 <= '0';
			b2 <= '0';
			b3 <= '1';
			b4 <= '0';
			b5 <= '0';
			b6 <= '0';
			elsif (rightMBs = "1011") then
			b0 <= '1';
			b1 <= '1';
			b2 <= '0';
			b3 <= '0';
			b4 <= '0';
			b5 <= '0';
			b6 <= '0';
			elsif (rightMBs = "1100") then
			b0 <= '0';
			b1 <= '1';
			b2 <= '1';
			b3 <= '0';
			b4 <= '0';
			b5 <= '0';
			b6 <= '1';
			elsif (rightMBs = "1101") then
			b0 <= '1';
			b1 <= '0';
			b2 <= '0';
			b3 <= '0';
			b4 <= '0';
			b5 <= '1';
			b6 <= '0';
			elsif (rightMBs = "1110") then
			b0 <= '0';
			b1 <= '1';
			b2 <= '1';
			b3 <= '0';
			b4 <= '0';
			b5 <= '0';
			b6 <= '0';
			elsif (rightMBs = "1111") then
			b0 <= '0';
			b1 <= '1';
			b2 <= '1';
			b3 <= '1';
			b4 <= '0';
			b5 <= '0';
			b6 <= '0';
		end if;
		
	end process;
	
	--for left display
	process (al_value) is
	begin
		if(leftMBs = "0000") then
			a0 <= '0';
			a1 <= '0';
			a2 <= '0';
			a3 <= '0';
			a4 <= '0';
			a5 <= '0';
			a6 <= '1';
		elsif (leftMBs = "0001") then
			a0 <= '1';
			a1 <= '0';
			a2 <= '0';
			a3 <= '1';
			a4 <= '1';
			a5 <= '1';
			a6 <= '1';
		elsif (leftMBs = "0010") then
			a0 <= '0';
			a1 <= '0';
			a2 <= '1';
			a3 <= '0';
			a4 <= '0';
			a5 <= '1';
			a6 <= '0';
		elsif (leftMBs = "0011") then
			a0 <= '0';
			a1 <= '0';
			a2 <= '0';
			a3 <= '0';
			a4 <= '1';
			a5 <= '1';
			a6 <= '0';
		elsif (leftMBs = "0100") then
			a0 <= '1';
			a1 <= '0';
			a2 <= '0';
			a3 <= '1';
			a4 <= '1';
			a5 <= '0';
			a6 <= '0';
		elsif (leftMBs = "0101") then
			a0 <= '0';
			a1 <= '1';
			a2 <= '0';
			a3 <= '0';
			a4 <= '1';
			a5 <= '0';
			a6 <= '0';
		elsif (leftMBs = "0110") then
			a0 <= '0';
			a1 <= '1';
			a2 <= '0';
			a3 <= '0';
			a4 <= '0';
			a5 <= '0';
			a6 <= '0';
		elsif (leftMBs = "0111") then
			a0 <= '0';
			a1 <= '0';
			a2 <= '0';
			a3 <= '1';
			a4 <= '1';
			a5 <= '1';
			a6 <= '1';
		elsif (leftMBs = "1000") then
			a0 <= '0';
			a1 <= '0';
			a2 <= '0';
			a3 <= '0';
			a4 <= '0';
			a5 <= '0';
			a6 <= '0';
		elsif (leftMBs = "1001") then
			a0 <= '0';
			a1 <= '0';
			a2 <= '0';
			a3 <= '1';
			a4 <= '1';
			a5 <= '0';
			a6 <= '0';
		elsif (leftMBs = "1010") then
			a0 <= '0';
			a1 <= '0';
			a2 <= '0';
			a3 <= '1';
			a4 <= '0';
			a5 <= '0';
			a6 <= '0';
		elsif (leftMBs = "1011") then
			a0 <= '1';
			a1 <= '1';
			a2 <= '0';
			a3 <= '0';
			a4 <= '0';
			a5 <= '0';
			a6 <= '0';
		elsif (leftMBs = "1100") then
			a0 <= '0';
			a1 <= '1';
			a2 <= '1';
			a3 <= '0';
			a4 <= '0';
			a5 <= '0';
			a6 <= '1';
		elsif (leftMBs = "1101") then
			a0 <= '1';
			a1 <= '0';
			a2 <= '0';
			a3 <= '0';
			a4 <= '0';
			a5 <= '1';
			a6 <= '0';
		elsif (leftMBs = "1110") then
			a0 <= '0';
			a1 <= '1';
			a2 <= '1';
			a3 <= '0';
			a4 <= '0';
			a5 <= '0';
			a6 <= '0';
		elsif (leftMBs = "1111") then
			a0 <= '0';
			a1 <= '1';
			a2 <= '1';
			a3 <= '1';
			a4 <= '0';
			a5 <= '0';
			a6 <= '0';
		end if;
		
	end process;

end rtl;
